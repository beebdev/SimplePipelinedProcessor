----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 29.03.2020 13:18:57
-- Design Name: 
-- Module Name: register_file - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity register_file is
    Port ( reset : in STD_LOGIC;
           clk : in STD_LOGIC;
           read_register_a : in STD_LOGIC_VECTOR (3 downto 0);
           read_register_b : in STD_LOGIC_VECTOR (3 downto 0);
           write_enable : in STD_LOGIC;
           write_register : in STD_LOGIC_VECTOR (3 downto 0);
           write_data : in STD_LOGIC_VECTOR (15 downto 0);
           read_data_a : out STD_LOGIC_VECTOR (15 downto 0);
           read_data_b : out STD_LOGIC_VECTOR (15 downto 0));
end register_file;

architecture Behavioral of register_file is

begin


end Behavioral;
